library verilog;
use verilog.vl_types.all;
entity Problem_2_vlg_vec_tst is
end Problem_2_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity DecoderDiagram_vlg_vec_tst is
end DecoderDiagram_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity ALU_1_vlg_vec_tst is
end ALU_1_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity FSMDiagram_vlg_vec_tst is
end FSMDiagram_vlg_vec_tst;
